module uwu

fn C.fgetc(&C.FILE) int
