module argser

pub struct Argser {
  ref &app.App
  args []string
}
